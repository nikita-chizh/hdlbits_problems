SELECTOR UNIQUE_CASE
UNIQUE_CASE FALSE
TEST_CASE LEADING_ONES