module top_module (
    input [4:0] a, b, c, d, e, f,
    output [7:0] w, x, y, z );
    wire [29:0] temp;
    assign temp = { a, b, c, d, e, f};
    assign {w, x, y, z} = {temp, 2'b11};

endmodule
