module top_module ( input a, input b, output out );
    mod_a mod_a_instance(a, b, out);
endmodule
